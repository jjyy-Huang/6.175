import Multiplexer::*;

// Full adder functions

function Bit#(1) fa_sum( Bit#(1) a, Bit#(1) b, Bit#(1) c_in );
    return xor1( xor1( a, b ), c_in );
endfunction

function Bit#(1) fa_carry( Bit#(1) a, Bit#(1) b, Bit#(1) c_in );
    return or1( and1( a, b ), and1( xor1( a, b ), c_in ) );
endfunction

// 4 Bit full adder

function Bit#(5) add4( Bit#(4) a, Bit#(4) b, Bit#(1) c_in );
    return 0;
endfunction

// Adder interface

interface Adder8;
    method ActionValue#( Bit#(9) ) sum( Bit#(8) a, Bit#(8) b, Bit#(1) c_in );
endinterface

// Adder modules

// RC = Ripple Carry
module mkRCAdder( Adder8 );
    method ActionValue#( Bit#(9) ) sum( Bit#(8) a, Bit#(8) b, Bit#(1) c_in );
        Bit#(5) lower_result = add4( a[3:0], b[3:0], c_in );
        Bit#(5) upper_result = add4( a[7:4], b[7:4], lower_result[4] );
        return { upper_result , lower_result[3:0] };
    endmethod
endmodule

// CS = Carry Select
module mkCSAdder( Adder8 );
    method ActionValue#( Bit#(9) ) sum( Bit#(8) a, Bit#(8) b, Bit#(1) c_in );
        return 0;
    endmethod
endmodule


// function Bit#(2) halfAdder(Bit#(1) aIn, Bit#(1) bIn);
//   let sOut = aIn ^ bIn;
//   let cOut = aIn & bIn;
//   return {cOut, sOut};
// endfunction

// function Bit#(2) fullAdder(Bit#(1) aIn, Bit#(1) bIn, Bit#(1) cIn);
//   let ab = halfAdder(aIn, bIn);
//   let abc = halfAdder(ab[0], cIn);
//   let sOut = abc[0];
//   let cOut = abc[1] | ab[1];
//   return {cOut, sOut};

// endfunction

// function Bit#(TAdd#(width, 1)) ripplerAdderN(Bit#(width) aIn, Bit#(width) bIn, Bit#(1) cIn);
//   Bit#(width) sOut;
//   Bit#(TAdd#(width, 1)) carry;
//   carry[0] = cIn;
//   let widthValue = valueOf(width);
//   for( Integer idx = 0; idx < widthValue; idx = idx + 1) begin
//     let cs = fullAdder(aIn[idx], bIn[idx], carry[idx]);
//     sOut[idx] = cs[0];
//     carry[idx + 1] = cs[1];
//   end
//   return {carry[widthValue], sOut};
// endfunction

// function Bit#(5) add4( Bit#(4) a, Bit#(4) b, Bit#(1) c_in );
//     Bit#(4) s; Bit#(5) c = 0; c[0] = c_in;
//     for(Integer i = 0; i < 4; i = i + 1) begin
//         s[i] = fa_sum(a[i], b[i], c[i]);
//         c[i+1] = fa_carry(a[i], b[i], c[i]);
//     end
//     return { c[4], s };
// endfunction
